module test2;
 logic [3:0] a1;
 logic red1,green1,blue1;

task1 aa_b (
   .a(a1),
   .red(red1),
   .green(green1),
   .blue(blue1)

 );

 initial begin
    
    a1[3] = 0 ; a1[2] = 0; a1[1] = 0; a1[0] = 0;
    #10;
    a1[3] = 0; a1[2] = 0; a1[1] = 0; a1[0]=1;
    #10;
    a1[3] = 0; a1[2] = 0; a1[1] = 1; a1[0]=0;
    #10;
    a1[3] = 0; a1[2] = 0; a1[1] = 1; a1[0]=1;
    #10;
    a1[3] = 0; a1[2] = 1; a1[1] = 0; a1[0]=0;
    #10;
    a1[3] = 0; a1[2] = 1; a1[1] = 0; a1[0]=1;
    #10;
    a1[3] = 0; a1[2] = 1; a1[1] = 1; a1[0]=0;
    #10;
    a1[3] = 0; a1[2] = 1; a1[1] = 1; a1[0]=1;
    #10;
    a1[3] = 1; a1[2] = 0; a1[1] = 0; a1[0]=0;
    #10;
    a1[3] = 1; a1[2] = 0; a1[1] = 0; a1[0]=1;
    #10;
    a1[3] = 1; a1[2] = 0; a1[1] = 1; a1[0]=0;
    #10;
    a1[3] = 1; a1[2] = 0; a1[1] = 1; a1[0]=1;
    #10;
    a1[3] = 1; a1[2] = 1; a1[1] = 0; a1[0]=0;
    #10;
    a1[3] = 1; a1[2] = 1; a1[1] = 0; a1[0]=1;
    #10;
    a1[3] = 1; a1[2] = 1; a1[1] = 1; a1[0]=0;
    #10;
    a1[3] = 1; a1[2] = 1; a1[1] = 1; a1[0]=1;
    #10;
    $stop;
 end

 endmodule